module and_g(input logic a,input logic b,output logic c);

assign c=a&b;
endmodule

